// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

`define ETHERNET_XXVGMII_CLOCK                      1280
`define ETHERNET_SERIAL_CAUI_25G_CLOCK              (19.3939)
`define ETHERNET_XXVSBI_CLOCK                       (620.608/2)
`define ETHERNET_REFERENCE_CLOCK                    50 
`define ETHERNET_GMII_CLOCK                         4000
`define ETHERNET_SERIAL_BASER_CLOCK                 (96.97/2.0) 
`define ETHERNET_SERIAL_BASE4X_CLOCK                160
`define ETHERNET_SERIAL_BASEX_CLOCK                 400
`define ETHERNET_GMII_CLOCK                         4000
`define ETHERNET_25MHZ_CLOCK                        20000
`define ETHERNET_2PT5_MHZ_CLOCK                     200000
`define ETHERNET_SGMII_CLOCK                        80
`define ETHERNET_QSGMII_CLOCK                       100
`define ETHERNET_TBI_CLOCK                          4000
`define ETHERNET_XLGMII_CLOCK                       800
`define ETHERNET_XXGMII_CLOCK                       1600
`define ETHERNET_CGMII_CLOCK                        320
`define ETHERNET_CGMII_MIMIC_DUT_CLOCK              160
`define ETHERNET_XLGMII_MIMIC_DUT_CLOCK             400
`define ETHERNET_XGMII_CLOCK                        3200
`define ETHERNET_FBI_CLOCK                          1600
`define ETHERNET_SERIAL_CLOCK_BASEX                 40
`define ETHERNET_XSBI_CLOCK                         (1551.52/2.0)
`define ETHERNET_VSBI_CLOCK                         1551.52
`define ETHERNET_VSBI_CLOCK_CAUI_25x4_64B_PARALLEL  (3103.03/2.0)
`define ETHERNET_CAUI_64B_PARALLEL_CLOCK            (2482.424/2)   
`define ETHERNET_REFERENCE_CLOCK                    50 
`define ETHERNET_KR4_FEC_66_CLOCK                   1280
`define ETHERNET_KR4_FEC_40_CLOCK                   775.757576
`define ETHERNET_ROUND_TRIP_TIME                    4000
`define ETHERNET_RMII_CLOCK                         10000
`define ETHERNET_GMII_RMII_CLOCK                    40000
`define ETHERNET_MDIO_CLOCK                         200
`define ETHERNET_PTP_SYS_CLOCK                      500000
`define ETHERNET_XXVGMII_CLOCK                      1280
`define ETHERNET_LGMII_CLOCK                        640
`define ETHERNET_XXVSBI_CLOCK                       (620.608/2)
`define ETHERNET_LSBI_CLOCK                         (620.608)
`define ETHERNET_SERIAL_12pt5G_CLOCK                (38.788)
`define ETHERNET_SERIAL_CD_CLOCK                    18.824
`define ETHERNET_SERIAL_50G_CLOCK                   9.412
`define ETHERNET_CDMII_CLOCK                        80
`define ETHERNET_CCMII_CLOCK                        160
`define ETHERNET_CDXBI_CLOCK                        (376.48/2)
