pmci_csr_test
pmci_qsfp_telemetry_test
pmci_multi_master_test
pmci_mailbox_test
pmci_ro_mailbox_test
pmci_vdm_tx_rx_lpbk_test
pmci_vdm_mctp_mmio_b2b_test
pmci_rd_default_value_test
pmci_vdm_tlp_error_scenario_test
pmci_vdm_b2b_drop_err_scenario_test
pmci_vdm_len_err_scenario_test
pmci_vdm_multipkt_error_scenario_test
pmci_vdm_multipkt_tlp_err_test
pmci_vdm_tx_rx_all_toggle_test
pmci_vdm_tx_rx_all_random_lpbk_test
