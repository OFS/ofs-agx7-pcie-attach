// Copyright (C) 2021 Intel Corporation.
// SPDX-License-Identifier: MIT

//
// Description
//-----------------------------------------------------------------------------
//
// This package defines the FIM clk for BASE_X16_ADP
//
//----------------------------------------------------------------------------

`ifndef __OFS_AXI_FIM_CLK_PKG_SV__
`define __OFS_AXI_FIM_CLK_PKG_SV__

package ofs_axi_fim_clk_pkg;

localparam AXI_FIM_CLK_HZ = 400000000; //400MHz

endpackage

`endif // __OFS_AXI_FIM_CLK_PKG_SV__
