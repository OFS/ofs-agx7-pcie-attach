//Copyright (C) 2021 Intel Corporation
//SPDX-License-Identifier: MIT
`ifndef TX_TEST_PKG_100G_200G_SVH
`define TX_TEST_PKG_100G_200G_SVH

//package test_pkg;
//    import uvm_pkg::*;
//    `include "uvm_macros.svh"

    `include "base_test.svh"
    `include "he_hssi_tx_lpbk_P0_test.svh"
    `include "he_hssi_tx_lpbk_P1_test.svh"

    //endpackage : test_pkg

`endif // TX_TEST_PKG_100G_200G_SVH
