//Copyright (C) 2021 Intel Corporation
//SPDX-License-Identifier: MIT
`ifndef TX_TEST_PKG_SVH
`define TX_TEST_PKG_SVH

//package test_pkg;
//    import uvm_pkg::*;
//    `include "uvm_macros.svh"

    `include "base_test.svh"
    `include "he_hssi_csr_test.svh"
    `include "he_hssi_axis_rx_lpbk_test.svh"
    `include "he_hssi_tx_lpbk_P0_test.svh"
    `include "he_hssi_tx_lpbk_P1_test.svh"
    `include "he_hssi_tx_lpbk_P2_test.svh"
    `include "he_hssi_tx_lpbk_P3_test.svh"
    `include "he_hssi_tx_lpbk_P4_test.svh"
    `include "he_hssi_tx_lpbk_P5_test.svh"
    `include "he_hssi_tx_lpbk_P6_test.svh"
    `include "he_hssi_tx_lpbk_P7_test.svh"
    `include "he_hssi_tx_err_L0_test.svh"
    `include "he_hssi_tx_err_L1_test.svh"
    `include "he_hssi_tx_err_L2_test.svh"
    `include "he_hssi_tx_err_L3_test.svh"
    `include "he_hssi_tx_err_L4_test.svh"
    `include "he_hssi_tx_err_L5_test.svh"
    `include "he_hssi_tx_err_L6_test.svh"
    `include "he_hssi_tx_err_L7_test.svh"

    //endpackage : test_pkg

`endif // TX_TEST_PKG_SVH
