//Copyright (C) 2021 Intel Corporation
//SPDX-License-Identifier: MIT
`ifndef RX_TEST_PKG_100G_SVH
`define RX_TEST_PKG_100G_SVH

//package test_pkg;
//    import uvm_pkg::*;
//    `include "uvm_macros.svh"
   `include "base_test.svh"
   `include "he_hssi_rx_lpbk_100G_test.svh"
`endif // RX_TEST_PKG_100G_SVH
