// Copyright (C) 2021 Intel Corporation
// SPDX-License-Identifier: MIT

// i2c_bfm.v

// Generated using ACDS version 20.1 177

`timescale 1 ps / 1 ps
module i2c_bfm (
		input  wire        clk,           //         clock.clk
		output wire [31:0] address,       // avalon_master.address
		output wire        read,          //              .read
		input  wire [31:0] readdata,      //              .readdata
		input  wire        readdatavalid, //              .readdatavalid
		input  wire        waitrequest,   //              .waitrequest
		output wire        write,         //              .write
		output wire [3:0]  byteenable,    //              .byteenable
		output wire [31:0] writedata,     //              .writedata
		input  wire        rst_n,         //         reset.reset_n
		input  wire        i2c_data_in,   //   conduit_end.conduit_data_in
		input  wire        i2c_clk_in,    //              .conduit_clk_in
		output wire        i2c_data_oe,   //              .conduit_data_oe
		output wire        i2c_clk_oe     //              .conduit_clk_oe
	);

	altera_i2cslave_to_avlmm_bridge #(
		.I2C_SLAVE_ADDRESS (7'b1010000),
		.BYTE_ADDRESSING   (1),
		.ADDRESS_STEALING  (0),
		.READ_ONLY         (0)
	) i2cslave_to_avlmm_bridge_0 (
		.clk           (clk),           //   input,   width = 1,         clock.clk
		.address       (address),       //  output,  width = 32, avalon_master.address
		.read          (read),          //  output,   width = 1,              .read
		.readdata      (readdata),      //   input,  width = 32,              .readdata
		.readdatavalid (readdatavalid), //   input,   width = 1,              .readdatavalid
		.waitrequest   (waitrequest),   //   input,   width = 1,              .waitrequest
		.write         (write),         //  output,   width = 1,              .write
		.byteenable    (byteenable),    //  output,   width = 4,              .byteenable
		.writedata     (writedata),     //  output,  width = 32,              .writedata
		.rst_n         (rst_n),         //   input,   width = 1,         reset.reset_n
		.i2c_data_in   (i2c_data_in),   //   input,   width = 1,   conduit_end.conduit_data_in
		.i2c_clk_in    (i2c_clk_in),    //   input,   width = 1,              .conduit_clk_in
		.i2c_data_oe   (i2c_data_oe),   //  output,   width = 1,              .conduit_data_oe
		.i2c_clk_oe    (i2c_clk_oe)     //  output,   width = 1,              .conduit_clk_oe
	);

endmodule
